--  This is a top level module for our system
-- *Configuration can be changed from this file